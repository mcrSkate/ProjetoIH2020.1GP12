module inst_concatener (
    input wire [15:0] Instr15_0;
    input wire [4:0] Instr20_16;
);
    
endmodule