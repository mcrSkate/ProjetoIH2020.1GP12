module div (
    input wire [31:0] regA_out;
    input wire [31:0] regB_out;
    input wire clock;
    input wire reset;
    input wire divControl;
    output wire zeroDiv
);
    
endmodule